interface interfaz (input clk);
  logic [2:0] r_mode;
  logic [32:0] fp_X;
  logic [32:0] fp_Y;
  logic [32:0] fp_Z;
  logic ovrf;
  logic udrf;
endinterface